module logic_gates(input a,b,output c);
and and1(c,a,b);
endmodule

